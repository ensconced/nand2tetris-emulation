module not_gate (input in,
                output out);
    nand_gate NANDA (in, in, out);
endmodule
